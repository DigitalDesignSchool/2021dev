`include "multi_memory.sv"
