

`include "fifo_w8.sv"

